module clock (
    output clk
);

    
    
endmodule